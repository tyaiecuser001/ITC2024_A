`timescale 1ns/100ps
module testbench;

reg iCLK,RST_n,rx,tx_en;

wire [7:0] LED;
wire tx,Server_wifi_txd;

TOP UART_Server(
			.iCLK(iCLK),
			.RST_n(RST_n),
			.tx_en(tx_en),
			.rx(rx),
			.tx(tx),
			.LED(LED),
			.Server_wifi_txd(Server_wifi_txd)
			);

initial
	begin
		iCLK <= 1'd1;
		RST_n <= 1'd0;
		rx <= 1'd1;
		tx_en <= 1'd0;
	end
	
initial
forever
	#10 iCLK = ~iCLK;
	

initial
	begin
		#60000 RST_n <= 1'd1; tx_en <= 1'd1;
		#1250000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#1500000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#3500000		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#2000000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#2000000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#4000000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#2000000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#2000000 		rx <= 1'd0;//43
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4e
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4e
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//45
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//43
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//54
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		
		#6000000 		rx <= 1'd0;//33h
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#6000000 $finish;
	end

endmodule
