`timescale 1ns/100ps
module testbench;

reg iCLK,RST_n,rx,select;
reg [3:0] SW;

wire Client_wifi_txd;


TOP TOP_u1(
			.iCLK(iCLK),
			.RST_n(RST_n),
			.select(select),
			.rx(rx),
			.SW(SW),
			.tx(tx),
			.Client_wifi_txd(Client_wifi_txd)
			);
			
			
initial
	begin
		iCLK <= 1'd1;
		RST_n <=1'd0;
		rx <= 1'd1;
		select <= 1'd1;
		SW <= 4'd1;
	end
	
initial
forever
	#10 iCLK = ~iCLK;
initial
	begin
		#120000 RST_n <= 1'd1;
		#1250000 		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#3000000		rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#3500000 	rx <= 1'd0;//4f   5
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1; 
		
		#2000000		SW <= 4'd3;
		#8660			select <= 1'd0;
		#125000			select <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;

#2000000		SW <= 4'd0;
		#8660			select <= 1'd0;
		#125000			select <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#2000000 	rx <= 1'd0;//4f
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//4b
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0d
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;//0a
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd0;
		#8660 		rx <= 1'd1;		
		
		#6000000 $finish;
	end
endmodule
